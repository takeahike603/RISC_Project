module ajc_8bit_const_unit_v (Func_Sel, Const_Result, Const_CNVZ);
//----------------------------------------------------------------------------------
// Input and output ports declarations
//----------------------------------------------------------------------------------
	input [1:0] Func_Sel;
	output [7:0] Const_Result; 
	output [3:0] Const_CNVZ;
//----------------------------------------------------------------------------------
// The const_mux instance
//----------------------------------------------------------------------------------
	ajc_nbit_4to1mux_v #8	const_mux
		(8'b11111111, 8'b10101010, 8'b01010101, 8'b00000000, Func_Sel[1:0], Const_Result);
//----------------------------------------------------------------------------------
	assign Const_CNVZ = {1'b0, Const_Result[3], 1'b0, ~| Const_Result};
//----------------------------------------------------------------------------------
endmodule
